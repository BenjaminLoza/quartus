library verilog;
use verilog.vl_types.all;
entity ParteF_vlg_vec_tst is
end ParteF_vlg_vec_tst;
