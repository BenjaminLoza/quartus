library verilog;
use verilog.vl_types.all;
entity ParteB is
    port(
        D               : in     vl_logic;
        CL              : in     vl_logic;
        Q               : out    vl_logic
    );
end ParteB;
