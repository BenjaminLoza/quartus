library verilog;
use verilog.vl_types.all;
entity ParteDstate_vlg_vec_tst is
end ParteDstate_vlg_vec_tst;
