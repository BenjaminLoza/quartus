-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- PROGRAM		"Quartus II 64-Bit"
-- VERSION		"Version 13.1.0 Build 162 10/23/2013 SJ Web Edition"
-- CREATED		"Wed Nov 06 20:26:37 2024"

LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

ENTITY dir IS 
	PORT
	(
		sda :  IN  STD_LOGIC;
		hdi :  IN  STD_LOGIC;
		rs :  IN  STD_LOGIC;
		clk :  IN  STD_LOGIC;
		fdi :  OUT  STD_LOGIC;
		soy :  OUT  STD_LOGIC
	);
END dir;

ARCHITECTURE bdf_type OF dir IS 

SIGNAL	SYNTHESIZED_WIRE_0 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_43 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_44 :  STD_LOGIC;
SIGNAL	DFF_inst9 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_45 :  STD_LOGIC;
SIGNAL	DFF_inst10 :  STD_LOGIC;
SIGNAL	DFF_inst11 :  STD_LOGIC;
SIGNAL	DFF_inst12 :  STD_LOGIC;
SIGNAL	DFF_inst13 :  STD_LOGIC;
SIGNAL	DFF_inst14 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_46 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_47 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_48 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_49 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_50 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_51 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_52 :  STD_LOGIC;
SIGNAL	DFF_inst8 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_22 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_23 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_24 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_25 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_26 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_27 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_28 :  STD_LOGIC;


BEGIN 
fdi <= SYNTHESIZED_WIRE_43;
SYNTHESIZED_WIRE_45 <= '1';
SYNTHESIZED_WIRE_47 <= '1';



SYNTHESIZED_WIRE_44 <= hdi AND SYNTHESIZED_WIRE_0 AND clk;


SYNTHESIZED_WIRE_0 <= NOT(SYNTHESIZED_WIRE_43);



PROCESS(SYNTHESIZED_WIRE_44,rs,SYNTHESIZED_WIRE_45)
BEGIN
IF (rs = '0') THEN
	DFF_inst10 <= '0';
ELSIF (SYNTHESIZED_WIRE_45 = '0') THEN
	DFF_inst10 <= '1';
ELSIF (RISING_EDGE(SYNTHESIZED_WIRE_44)) THEN
	DFF_inst10 <= DFF_inst9;
END IF;
END PROCESS;


PROCESS(SYNTHESIZED_WIRE_44,rs,SYNTHESIZED_WIRE_45)
BEGIN
IF (rs = '0') THEN
	DFF_inst11 <= '0';
ELSIF (SYNTHESIZED_WIRE_45 = '0') THEN
	DFF_inst11 <= '1';
ELSIF (RISING_EDGE(SYNTHESIZED_WIRE_44)) THEN
	DFF_inst11 <= DFF_inst10;
END IF;
END PROCESS;


PROCESS(SYNTHESIZED_WIRE_44,rs,SYNTHESIZED_WIRE_45)
BEGIN
IF (rs = '0') THEN
	DFF_inst12 <= '0';
ELSIF (SYNTHESIZED_WIRE_45 = '0') THEN
	DFF_inst12 <= '1';
ELSIF (RISING_EDGE(SYNTHESIZED_WIRE_44)) THEN
	DFF_inst12 <= DFF_inst11;
END IF;
END PROCESS;


PROCESS(SYNTHESIZED_WIRE_44,rs,SYNTHESIZED_WIRE_45)
BEGIN
IF (rs = '0') THEN
	DFF_inst13 <= '0';
ELSIF (SYNTHESIZED_WIRE_45 = '0') THEN
	DFF_inst13 <= '1';
ELSIF (RISING_EDGE(SYNTHESIZED_WIRE_44)) THEN
	DFF_inst13 <= DFF_inst12;
END IF;
END PROCESS;


PROCESS(SYNTHESIZED_WIRE_44,rs,SYNTHESIZED_WIRE_45)
BEGIN
IF (rs = '0') THEN
	DFF_inst14 <= '0';
ELSIF (SYNTHESIZED_WIRE_45 = '0') THEN
	DFF_inst14 <= '1';
ELSIF (RISING_EDGE(SYNTHESIZED_WIRE_44)) THEN
	DFF_inst14 <= DFF_inst13;
END IF;
END PROCESS;


PROCESS(SYNTHESIZED_WIRE_44,rs,SYNTHESIZED_WIRE_45)
BEGIN
IF (rs = '0') THEN
	SYNTHESIZED_WIRE_43 <= '0';
ELSIF (SYNTHESIZED_WIRE_45 = '0') THEN
	SYNTHESIZED_WIRE_43 <= '1';
ELSIF (RISING_EDGE(SYNTHESIZED_WIRE_44)) THEN
	SYNTHESIZED_WIRE_43 <= DFF_inst14;
END IF;
END PROCESS;



SYNTHESIZED_WIRE_27 <= SYNTHESIZED_WIRE_46 AND SYNTHESIZED_WIRE_47;


SYNTHESIZED_WIRE_25 <= SYNTHESIZED_WIRE_48 AND SYNTHESIZED_WIRE_47;


SYNTHESIZED_WIRE_26 <= SYNTHESIZED_WIRE_49 AND SYNTHESIZED_WIRE_47;


PROCESS(SYNTHESIZED_WIRE_44,rs,SYNTHESIZED_WIRE_45)
BEGIN
IF (rs = '0') THEN
	SYNTHESIZED_WIRE_46 <= '0';
ELSIF (SYNTHESIZED_WIRE_45 = '0') THEN
	SYNTHESIZED_WIRE_46 <= '1';
ELSIF (RISING_EDGE(SYNTHESIZED_WIRE_44)) THEN
	SYNTHESIZED_WIRE_46 <= sda;
END IF;
END PROCESS;


SYNTHESIZED_WIRE_28 <= SYNTHESIZED_WIRE_50 AND SYNTHESIZED_WIRE_47;


SYNTHESIZED_WIRE_24 <= SYNTHESIZED_WIRE_51 AND SYNTHESIZED_WIRE_47;


SYNTHESIZED_WIRE_22 <= SYNTHESIZED_WIRE_52 AND SYNTHESIZED_WIRE_47;


SYNTHESIZED_WIRE_23 <= DFF_inst8 AND SYNTHESIZED_WIRE_47;



soy <= SYNTHESIZED_WIRE_43 AND SYNTHESIZED_WIRE_22 AND SYNTHESIZED_WIRE_23 AND SYNTHESIZED_WIRE_24 AND SYNTHESIZED_WIRE_25 AND SYNTHESIZED_WIRE_26 AND SYNTHESIZED_WIRE_27 AND SYNTHESIZED_WIRE_28;


PROCESS(SYNTHESIZED_WIRE_44,rs)
BEGIN
IF (rs = '0') THEN
	SYNTHESIZED_WIRE_48 <= '0';
ELSIF (RISING_EDGE(SYNTHESIZED_WIRE_44)) THEN
	SYNTHESIZED_WIRE_48 <= SYNTHESIZED_WIRE_46;
END IF;
END PROCESS;


PROCESS(SYNTHESIZED_WIRE_44,rs,SYNTHESIZED_WIRE_45)
BEGIN
IF (rs = '0') THEN
	SYNTHESIZED_WIRE_49 <= '0';
ELSIF (SYNTHESIZED_WIRE_45 = '0') THEN
	SYNTHESIZED_WIRE_49 <= '1';
ELSIF (RISING_EDGE(SYNTHESIZED_WIRE_44)) THEN
	SYNTHESIZED_WIRE_49 <= SYNTHESIZED_WIRE_48;
END IF;
END PROCESS;


PROCESS(SYNTHESIZED_WIRE_44,rs,SYNTHESIZED_WIRE_45)
BEGIN
IF (rs = '0') THEN
	SYNTHESIZED_WIRE_50 <= '0';
ELSIF (SYNTHESIZED_WIRE_45 = '0') THEN
	SYNTHESIZED_WIRE_50 <= '1';
ELSIF (RISING_EDGE(SYNTHESIZED_WIRE_44)) THEN
	SYNTHESIZED_WIRE_50 <= SYNTHESIZED_WIRE_49;
END IF;
END PROCESS;


PROCESS(SYNTHESIZED_WIRE_44,rs,SYNTHESIZED_WIRE_45)
BEGIN
IF (rs = '0') THEN
	SYNTHESIZED_WIRE_51 <= '0';
ELSIF (SYNTHESIZED_WIRE_45 = '0') THEN
	SYNTHESIZED_WIRE_51 <= '1';
ELSIF (RISING_EDGE(SYNTHESIZED_WIRE_44)) THEN
	SYNTHESIZED_WIRE_51 <= SYNTHESIZED_WIRE_50;
END IF;
END PROCESS;


PROCESS(SYNTHESIZED_WIRE_44,rs,SYNTHESIZED_WIRE_45)
BEGIN
IF (rs = '0') THEN
	SYNTHESIZED_WIRE_52 <= '0';
ELSIF (SYNTHESIZED_WIRE_45 = '0') THEN
	SYNTHESIZED_WIRE_52 <= '1';
ELSIF (RISING_EDGE(SYNTHESIZED_WIRE_44)) THEN
	SYNTHESIZED_WIRE_52 <= SYNTHESIZED_WIRE_51;
END IF;
END PROCESS;


PROCESS(SYNTHESIZED_WIRE_44,rs,SYNTHESIZED_WIRE_45)
BEGIN
IF (rs = '0') THEN
	DFF_inst8 <= '0';
ELSIF (SYNTHESIZED_WIRE_45 = '0') THEN
	DFF_inst8 <= '1';
ELSIF (RISING_EDGE(SYNTHESIZED_WIRE_44)) THEN
	DFF_inst8 <= SYNTHESIZED_WIRE_52;
END IF;
END PROCESS;


PROCESS(SYNTHESIZED_WIRE_44,rs,SYNTHESIZED_WIRE_45)
BEGIN
IF (rs = '0') THEN
	DFF_inst9 <= '0';
ELSIF (SYNTHESIZED_WIRE_45 = '0') THEN
	DFF_inst9 <= '1';
ELSIF (RISING_EDGE(SYNTHESIZED_WIRE_44)) THEN
	DFF_inst9 <= SYNTHESIZED_WIRE_45;
END IF;
END PROCESS;


END bdf_type;