library ieee;
use ieee.std_logic_1164.all;

entity ParteB is
	Port (
		D,CL: in std_logic;
		Q: out std_logic);
		end;
		
architecture behaviour of ParteB is
begin

end; 