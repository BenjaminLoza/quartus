library verilog;
use verilog.vl_types.all;
entity ParteB_vlg_vec_tst is
end ParteB_vlg_vec_tst;
